module circuito_autenticacao(a,b,c,d,e,f)




endmodule 