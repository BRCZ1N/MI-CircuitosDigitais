module circuito_comparador_funcionalidade(a,b,c,d,e,f)




endmodule 