module decodificador_7Seg(A,B,C);

	input A, B, C;


endmodule 