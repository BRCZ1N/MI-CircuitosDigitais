module circuito_codificador_autenticacao(a,b,c,d,e,f)




endmodule 