module decodificador_matriz(a,b,c,d,e,f)




endmodule 