module decodificador_matriz(A,B,C,MLED0,MLED1,LED2,LED3,LED4,LED5,LED6,LED7);

	input A, B, C;
	output MLED0,MLED1,LED2,LED3,LED4,LED5,LED6,LED7;
	wire NA = !A, NB = !B, NC = !C
	
	

endmodule 