module decodificador_7Seg(a,b,c,d,e,f)




endmodule 