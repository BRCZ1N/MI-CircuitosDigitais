module decodificador_leds(A,B,C);

	input A, B, C;


endmodule 