module circuito_seletor_saidas(a,b,c,d,e,f)




endmodule 