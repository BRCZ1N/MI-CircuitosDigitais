module circuito_seletor_7seg(A,B,C);

	input A, B, C;


endmodule 