module PBL_1(a,b,c,d,e,f)




endmodule 