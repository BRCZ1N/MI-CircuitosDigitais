module pbl(A,B,C);
	
	input A, B, C;



endmodule 