module circuito_7seg_f2(a,b,c,d,e,f)




endmodule 