module circuito_seletor_7seg(a,b,c,d,e,f)




endmodule 