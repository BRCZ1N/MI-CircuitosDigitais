module decodificador_matriz(A,B,C);

	input A, B, C;
	

endmodule 