module circuito_comparador_funcionalidade(A,B,C);	

	input A, B, C;


endmodule 