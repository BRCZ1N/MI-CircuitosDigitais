module circuito_comparador_autenticacao(A,B,C);

	input A, B, C;


endmodule 