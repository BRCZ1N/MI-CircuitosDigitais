module seletor_terminais(A,B,C);

	input A, B, C;


endmodule 