module mux2_1(A,B,C);

	input A, B, C;


endmodule 