module seletor_terminais(a,b,c,d,e,f)




endmodule 