module pbl(HH0,HH1,HH2,HH3,B3,B2,HH4,HH5,HH6,HH7,B1,B0,LED0,LED1,LED2,LED3,LED4,LED5,LED6,MLED0,MLED1,MLED2,MLED3,MLED4,MLED5,MLED6,MLED7,SEGA,SEGB,SEGC,SEGD,SEGE,SEGF,SEGG,SEGDP);
	
	input HH0,HH1,HH2,HH3,B3,B2,HH4,HH5,HH6,HH7,B1,B0;
	output LED0,LED1,LED2,LED3,LED4,LED5,LED6,MLED0,MLED1,MLED2,MLED3,MLED4,MLED5,MLED6,MLED7,SEGA,SEGB,SEGC,SEGD,SEGE,SEGF,SEGG,SEGDP;

endmodule 