module circuito_7seg_f2(A,B,C);

	input A, B, C;


endmodule 