module pbl(a,b,c,d,e,f)




endmodule 